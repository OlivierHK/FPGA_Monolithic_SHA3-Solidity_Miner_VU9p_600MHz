--------------------------------------------------------------------------------
-- PROJECT: ALTO FPGA Miner. SHA3-Solidity Flavor on Virtex ULTRAScale XCVU9P
--------------------------------------------------------------------------------
-- AUTHORS: Olivier FAURIE <olivier.faurie.hk@gmail.com>
-- LICENSE: 
-- WEBSITE: https://github.com/olivierHK
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.MATH_REAL.ALL;

Library UNISIM;
use UNISIM.vcomponents.all;

library work;
use work.MyPackage.all;



entity ROM_DRP_CLK_MODULE is
    Port ( 
    i_ROM_clk  : in  std_logic;
    i_ROM_en   : in  std_logic;
    i_ROM_addr : in  std_logic_vector(11 downto 0);
    o_ROM_data : out std_logic_vector(23 downto 0) 
    );
end entity;
------------------------------------------------------------------


architecture ROM_DRP_CLK_MODULE_arch of ROM_DRP_CLK_MODULE is

    type rom_type is array (0 to 4095) of std_logic_vector(23 downto 0); 
    
    signal ROM : rom_type := (  X"14179e",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081186",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081186",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416dc",  X"150080",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081186",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1415d7",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081186",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141820",  X"150000",  X"160104",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081104",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141659",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081186",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169a",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081186",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c4",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081104",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081105",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14175d",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081104",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179e",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081104",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417df",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081104",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141820",  X"150000",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081104",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416dc",  X"150080",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081104",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14165a",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081105",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141452",  X"150080",  X"160042",  X"4F9090",  X"4E9900",  X"27FFFF",  X"180113",  X"197c01",  X"1A7fe9",  X"081104",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c4",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141493",  X"150080",  X"160042",  X"4F9090",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081104",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14171d",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169a",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081104",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179e",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141515",  X"150080",  X"160082",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141556",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416dc",  X"150080",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179e",  X"150000",  X"160104",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1415d7",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1415d8",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141820",  X"150000",  X"160104",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141619",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141659",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14165a",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169a",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169b",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"0810c3",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c4",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416dc",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"160105",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14171d",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14175d",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14175e",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179e",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179f",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417df",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141820",  X"150000",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141820",  X"150000",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416dc",  X"150080",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416dc",  X"150080",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14165a",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1415d7",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141452",  X"150080",  X"160042",  X"4F9090",  X"4E9900",  X"27FFFF",  X"180113",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141452",  X"150080",  X"160042",  X"4F9090",  X"4E9900",  X"27FFFF",  X"180113",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c4",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c4",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141493",  X"150080",  X"160042",  X"4F9090",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141659",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14171d",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14171d",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169a",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169a",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081082",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179e",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416db",  X"150000",  X"160104",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141515",  X"150080",  X"160082",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141515",  X"150080",  X"160082",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141556",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14175d",  X"150000",  X"160104",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416dc",  X"150080",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416dc",  X"150080",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179e",  X"150000",  X"160104",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179e",  X"150000",  X"160104",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1415d7",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417df",  X"150000",  X"160104",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1415d8",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1415d8",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141820",  X"150000",  X"160104",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141820",  X"150000",  X"160104",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141619",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141411",  X"150080",  X"160082",  X"4F9090",  X"4E9900",  X"27FFFF",  X"18012c",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141659",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141659",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14165a",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14165a",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169a",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141452",  X"150080",  X"160082",  X"4F9090",  X"4E9900",  X"27FFFF",  X"180113",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169b",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169b",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081042",  X"090080",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c4",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c4",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416dc",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141493",  X"150080",  X"160082",  X"4F9090",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14171c",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14171c",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14171d",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14171d",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14175d",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1414d4",  X"150080",  X"160082",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14175e",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14175e",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179e",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179e",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179f",  X"150080",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141515",  X"150080",  X"160082",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417df",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417df",  X"150000",  X"1600c3",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1417e0",  X"150080",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141820",  X"150000",  X"1600c3",  X"4F1090",  X"4E9000",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141556",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141556",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141556",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416dc",  X"150080",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416dc",  X"150080",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1416dc",  X"150080",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141597",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141451",  X"150000",  X"160042",  X"4F9090",  X"4E9900",  X"27FFFF",  X"180113",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141451",  X"150000",  X"160042",  X"4F9090",  X"4E9900",  X"27FFFF",  X"180113",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1415d7",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1415d7",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141452",  X"150080",  X"160042",  X"4F9090",  X"4E9900",  X"27FFFF",  X"180113",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1415d8",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1415d8",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1415d8",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179e",  X"150000",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179e",  X"150000",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14179e",  X"150000",  X"160083",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141619",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141493",  X"150080",  X"160042",  X"4F9090",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141493",  X"150080",  X"160042",  X"4F9090",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141659",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141659",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"1414d3",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14165a",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14165a",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14165a",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169a",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169a",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169a",  X"150000",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"14169b",  X"150080",  X"160082",  X"4F0890",  X"4E9900",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000", 
                                X"141514",  X"150000",  X"160042",  X"4F0890",  X"4E9800",  X"27FFFF",  X"1800fa",  X"197c01",  X"1A7fe9",  X"081041",  X"090000",  X"000000",  X"000000",  X"000000",  X"000000",  X"000000" 


);  
    
    attribute rom_style : string;    
    attribute rom_style of ROM : signal is "block";
    
    begin   
    process(i_ROM_clk)  
        begin   
        if rising_edge(i_ROM_clk) then    
            if (i_ROM_en = '1') then    
                o_ROM_data <= ROM(conv_integer(i_ROM_addr));   
            end if;    
        end if;    
    end process; 
    
end architecture ROM_DRP_CLK_MODULE_arch;